library verilog;
use verilog.vl_types.all;
entity PRUEBA_vlg_vec_tst is
end PRUEBA_vlg_vec_tst;
