library verilog;
use verilog.vl_types.all;
entity VERIFICADOR_vlg_vec_tst is
end VERIFICADOR_vlg_vec_tst;
