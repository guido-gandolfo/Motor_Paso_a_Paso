library verilog;
use verilog.vl_types.all;
entity MOTORPAP_vlg_vec_tst is
end MOTORPAP_vlg_vec_tst;
