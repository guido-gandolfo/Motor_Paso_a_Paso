library verilog;
use verilog.vl_types.all;
entity FLIPFLOP_JK0_vlg_check_tst is
    port(
        SALIDA_Q0       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FLIPFLOP_JK0_vlg_check_tst;
