library verilog;
use verilog.vl_types.all;
entity FLIPFLOP_JK0_vlg_vec_tst is
end FLIPFLOP_JK0_vlg_vec_tst;
