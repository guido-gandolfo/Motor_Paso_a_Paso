library verilog;
use verilog.vl_types.all;
entity FLIPFLOP_JK1_vlg_check_tst is
    port(
        SALIDA_Q1       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FLIPFLOP_JK1_vlg_check_tst;
