library verilog;
use verilog.vl_types.all;
entity CONTROLADOR_COMPLETO_vlg_vec_tst is
end CONTROLADOR_COMPLETO_vlg_vec_tst;
