library verilog;
use verilog.vl_types.all;
entity FLIPFLOPJK2_vlg_check_tst is
    port(
        Q2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FLIPFLOPJK2_vlg_check_tst;
