library verilog;
use verilog.vl_types.all;
entity FLIPFLOPJK2_vlg_vec_tst is
end FLIPFLOPJK2_vlg_vec_tst;
