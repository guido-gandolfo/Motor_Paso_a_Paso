library verilog;
use verilog.vl_types.all;
entity FLIPFLOP_JK1_vlg_vec_tst is
end FLIPFLOP_JK1_vlg_vec_tst;
