library verilog;
use verilog.vl_types.all;
entity salidas_vlg_vec_tst is
end salidas_vlg_vec_tst;
