library verilog;
use verilog.vl_types.all;
entity MOTOR_vlg_vec_tst is
end MOTOR_vlg_vec_tst;
